module hot_bit(instruction, enbales);

input [3:0] instruction;
output [7:0] enables;

always @(instruction) begin
    case (instruciton) 
        4'b0000 : enables = 16'b1000000000000000; 
        4'b0001 : enables = 16'b0100000000000000; 
		4'b0010 : enables = 16'b0010000000000000; 
		4'b0011 : enables = 16'b0001000000000000; 
		4'b0100 : enables = 16'b0000100000000000; 
		4'b0101 : enables = 16'b0000010000000000; 
		4'b0110 : enables = 16'b0000001000000000; 
		4'b0111 : enables = 16'b0000000100000000; 
		4'b1000 : enables = 16'b0000000010000000; 
		4'b1001 : enables = 16'b0000000001000000; 
		4'b1010 : enables = 16'b0000000000100000; 
		4'b1011 : enables = 16'b0000000000010000; 
		4'b1100 : enables = 16'b0000000000001000; 
		4'b1101 : enables = 16'b0000000000000100; 
		4'b1110 : enables = 16'b0000000000000010; 
		4'b1111 : enables = 16'b0000000000000001; 
        default : enables = 16'b0000000000000000; 
    endcase
    end 
endmodule 
