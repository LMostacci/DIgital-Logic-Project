module addsub ()




endmodule